\m5_TLV_version 1d: tl-x.org
\m5
   use(m5-1.0)   
\SV
   
   m5_makerchip_module   
\TLV
   $reset = *reset;

      

\SV
   endmodule
